`define CMD_RDID 8'h9F
`define CMD_WRVECR 8'h61
`define CMD_WREN 8'h06
`define CMD_RFSR 8'h70
`define CMD_SE 8'hD8
`define CMD_BE 8'hC7
`define CMD_PP 8'h02

`define JEDEC_ID 8'h20

`define tPPmax 'd5 //ms
`define tBEmax 'd250_000 //ms
`define tSEmax 'd3_000 //ms
`define input_freq 'd40_000 //kHz
